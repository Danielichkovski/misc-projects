`timescale 1ns / 1ps
package my_testbench_pkg;
  import uvm_pkg::*;
  
  // The UVM sequence, transaction item, and driver are in these files:
  `include "my_transaction.svh"
  `include "my_scorboard.svh"
  `include "my_sequence.svh"
  `include "my_monitor.svh"
  `include "my_driver.svh"
  `include "my_agent.svh"
  `include "my_env.svh"
  `include "my_test.svh"
  

endpackage